module WolverineTest#(
                       parameter    NUM_MC_PORTS = 1,
                       parameter    RTNCTL_WIDTH = 32
                    )(
  input         clk,
  input         clkhx,
  input         clk2x,
  input         i_reset,
  input         disp_inst_vld,
  input  [4:0]  disp_inst,
  input  [17:0] disp_aeg_idx,
  input         disp_aeg_rd,
  input         disp_aeg_wr,
  input  [63:0] disp_aeg_wr_data,
  output [17:0] disp_aeg_cnt,
  output [15:0] disp_exception,
  output        disp_idle,
  output        disp_rtn_data_vld,
  output [63:0] disp_rtn_data,
  output        disp_stall,
  output        mc_rq_vld,
  output [31:0] mc_rq_rtnctl,
  output [63:0] mc_rq_data,
  output [47:0] mc_rq_vadr,
  output [1:0]  mc_rq_size,
  output [2:0]  mc_rq_cmd,
  output [3:0]  mc_rq_scmd,
  input         mc_rq_stall,
  input         mc_rs_vld,
  input  [2:0]  mc_rs_cmd,
  input  [3:0]  mc_rs_scmd,
  input  [63:0] mc_rs_data,
  input  [31:0] mc_rs_rtnctl,
  output        mc_rs_stall,
  output        mc_rq_flush,
  input         mc_rs_flush_cmplt,
  input         csr_wr_vld,
  input         csr_rd_vld,
  input  [15:0] csr_address,
  input  [63:0] csr_wr_data,
  output        csr_rd_ack,
  output [63:0] csr_rd_data,
  input  [3:0]  i_aeid
);
  WolverineShim top(
    .clock(clk),
    .reset(i_reset),
    .io_dispInstValid(disp_inst_vld),
    .io_dispInstData(disp_inst),
    .io_dispRegID(disp_aeg_idx),
    .io_dispRegRead(disp_aeg_rd),
    .io_dispRegWrite(disp_aeg_wr),
    .io_dispRegWrData(disp_aeg_wr_data),
    .io_dispAegCnt(disp_aeg_cnt),
    .io_dispException(disp_exception),
    .io_dispIdle(disp_idle),
    .io_dispRtnValid(disp_rtn_data_vld),
    .io_dispRtnData(disp_rtn_data),
    .io_dispStall(disp_stall),
    .io_mcReqValid(mc_rq_vld),
    .io_mcReqRtnCtl(mc_rq_rtnctl),
    .io_mcReqData(mc_rq_data),
    .io_mcReqAddr(mc_rq_vadr),
    .io_mcReqSize(mc_rq_size),
    .io_mcReqCmd(mc_rq_cmd),
    .io_mcReqSCmd(mc_rq_scmd),
    .io_mcReqStall(mc_rq_stall),
    .io_mcResValid(mc_rs_vld),
    .io_mcResCmd(mc_rs_cmd),
    .io_mcResSCmd(mc_rs_scmd),
    .io_mcResData(mc_rs_data),
    .io_mcResRtnCtl(mc_rs_rtnctl),
    .io_mcResStall(mc_rs_stall),
    .io_mcReqFlush(mc_rq_flush),
    .io_mcResFlushOK(mc_rs_flush_cmplt),
    .io_csrWrValid(csr_wr_vld),
    .io_csrRdValid(csr_rd_vld),
    .io_csrAddr(csr_address),
    .io_csrWrData(csr_wr_data),
    .io_csrReadAck(csr_rd_ack),
    .io_csrReadData(csr_rd_data),
    .io_aeid(i_aeid)
  );
endmodule